module dump();
    initial begin
        $dumpfile ("tt_um_tpu.vcd");
        $dumpvars (0, tt_um_tpu);
        #1;
    end
endmodule
