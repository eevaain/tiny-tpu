// HOW TO DIAGONALIZE INPUT DATA???

/*
- output only two elements at a time
- create a sort of program counter for each clock cycle? 
- program counter increments array value within whatever is loaded inside of this memory partition

*/

module input_setup(
    input [31:0] a11,
    input [31:0] a12, // inputs should be directly connected to 
    input [31:0] a21,
    input [31:0] a22,

    output [31:0] a_in1,
    output [31:0] a_in2
); 


always @(*) begin




    end


endmodule