`timescale 1ns / 1ns

/*  TODO: Figure out how to facilitate stream of data from computer to TPU 
^^ how can i move data from some memory partition from outside of my TPU, into my TPU. 
... Because at the moment I'm harcoding the weights and inputs.
*/

module tb_top_level_module;
  // Inputs
  reg clk;
  reg reset;
  reg [15:0] instruction;
  // Outputs
  wire [31:0] unified_mem [0:63];

  // Instantiate the top level module
  main uut (
    .clk(clk),
    .reset(reset),
    .instruction(instruction),
    .unified_mem(unified_mem)
  );

  // Clock generation
  always #5 clk = ~clk;

  // Initial block to initialize inputs and apply test vectors
  initial begin
    // Initialize inputs (registers outside the module)
    clk = 0;
    reset = 0;
    instruction = 0;

    // Apply reset (these are also registers outside the module)
    reset = 1;
    #10;
    reset = 0;
    #10;

    /// Load base address for weights (weights are in address 16 of WM)
    instruction = 16'b001_0000000001111;  // LOAD_ADDR 0x000F (16th address)
    #10;

    /// Load weights into systolic array
    instruction = 16'b010_0000000000000;  // LOAD_WEIGHT (Weights are transferred from weight memory into mmu)
    #10;

    /// Load base address for activation inputs (inputs start at address 30 of UB)
    instruction = 16'b001_0000000011110;  // LOAD_ADDR 0x001E (30th address)
    #10;

    /// Activation inputs are transferred from unified buffer to input setup unit
    instruction = 16'b011_0000000000000;  // LOAD_INPUT 
    #10;

    /// Convolutions begin within array. 
    instruction = 16'b100_0000000000000;  // COMPUTE (Compute starts, systolic operations are automated by here)

    #10; // now how can i get rid of this extra clock cycle?

    #10; // loads in a_in1 = 11; a_in2 = 0;
    #10; // loads in a_in1 = 12; a_in2 = 21;
    #10; // loads in a_in1 = 0; a_in2 = 22;

    #10; // mandatory empty input to allow partial sums to go into accumulator (i'm sure this one is mandatory)
    #10; // mandatory empty input to allow partial sums to go into accumulator (wait too sure about this one...)

    instruction = 16'b001_0000000000111;  // LOAD_ADDR 0x0007 (7th address)
    #10;

    // transfer accumulator product matrix rows into the unified buffer 
    instruction = 16'b101_0000000000000;  // STORE
    #10;

    // Monitor unified buffer
    $display("Unified Buffer at time %t:", $time);
    for (integer i = 0; i < 64; i = i + 1) begin
      $display("unified_mem[%0d] = %0d", i, unified_mem[i]);
    end

    // Finish the simulation
    $finish;
  end

endmodule
